Frequency vs Votage
.lib nom.lib
XA 0 2 3  4 5 2 7 4 555d
C 2 0 0.01u
C1 5 0 0.01U
RB 2 7 10K
RA 8 7 10K
VCC1 8 0 8
VCC 4 0 5V
RL 3 0 100K
.DC LIN VCC1 5 20 0.1
*1/((2.33* LOG10((3*V(8)-5)/(3* V(8)-10))*0.0002)+(0.000069))
.TRAN 20U 15M 0M 10U UIC
.PROBE
.END