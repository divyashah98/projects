
package simple_pkg;

    class my_class; 
        
        function new (string name);
            $display ("\nNAME is %s\n", name);
        endfunction
    endclass


endpackage
