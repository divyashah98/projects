// Defines parameters for various opcodes
localparam LDI  = 4'b0001;
localparam ADD  = 4'b0010;
localparam ADI  = 4'b0011;
localparam SUB  = 4'b0100;
localparam Mul  = 4'b0101;
localparam Div  = 4'b0110;
localparam INC  = 4'b0111;
localparam DEC  = 4'b1000;
localparam NOR  = 4'b1001;
localparam NAND = 4'b1010;
localparam XOR  = 4'b1011;
localparam COMP = 4'b1100;
localparam JMP  = 4'b1101;
localparam CMPJ = 4'b1110;
localparam NOP  = 4'b1111;
localparam HALT = 4'b0000;
