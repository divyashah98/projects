RC Phase Shift
.LIB EVAL.LIB
Xa 0 2 7 4 6 UA741
Vp 7 0 15
Vn 0 4 15
Rf 2 6 31K
Ra 2 1 1K
Ca 1 5 .01U
Rb 5 0 1K
Cb 5 9 .01U
Rc 9 0 1K
Cc 9 6 .01U
.TRAN 100U .5M
.PROBE
.END
