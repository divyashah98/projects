Band Reject Filter
.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
Ra 1 5 1K
Vp 7 0 15
Vn 0 4 15
Ca 5 0 2U
Rb 5 3 1K
Cb 1 8 1U
Cc 8 3 1U
Rc 8 6 0.5K
R2 6 2 0.9K
R1 2 0 1K
Vin 1 0 AC 100M
.AC DEC 20 10 10K
.PROBE
.END
