Input Offset Voltage R2 = 10K

.LIB EVAL.LIB
R1 0 2 100
R2 2 6 10K
V1 7 0 15
V2 0 4 15
X1 0 2 7 4 6 UA741
.END
