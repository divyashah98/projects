Schmitt Trigger Circuit(Hysteresis)
.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
R1 6 3 150K
R2 3 5 39K
Vref 5 0 0
Vin 1 0 pwl(0m 10 1m -10 2m 10)
Ron 2 1 31K
*Vin 1 0 AC 5 SIN(0 5 1K)
Rl 6 0 10K
Vp 7 0 15
Vn 0 4 15
.TRAN 100u 5M
.PROBE(V(6) V(3) V(1) V(5))
.END
