library verilog;
use verilog.vl_types.all;
entity pwm_tb is
end pwm_tb;
