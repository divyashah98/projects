Wein Bridge Oscillator
.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
Vp 7 0 15
Vn 0 4 15
Ri 2 0 1k
Rf 2 6 2.1K
C1 3 0 0.01U
R1 3 0 1K
C2 3 1 .01U
R2 1 6 1K
.TRAN 100U .2M
.PROBE
.END
