NON INVERTING AMPLIFIER

.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
V1 7 0 DC 15
V2 0 4 DC 15
Ra 2 0 1K
Rf 2 6 15K
Vs 3 0 AC 100M 90
Rl 6 0 10k
.AC LIN 10 10 100k
.PROBE
.END
