3.1 Open Loop Gain

.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
V0 3 0 DC 0
R4 2 3 10
R3 2 1 10K
R1 1 9 1.5K
RL 1 6 5.6K
V1 7 0 15
V2 0 4 15
Vs 9 0 DC 5
.DC Vs -5 5 .01
 
.PROBE
.END
