VOLTAGE FOLLOWER

.LIB EVAL.LIB
Xa 3 6 7 4 6 UA741
V1 0 4 15
V2 7 0 15
RL 6 0 10K
Vs 3 0 AC 100M 90
.AC LIN 100 100 1MEG
.PROBE
.END
