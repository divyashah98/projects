2.2 Bias And Offset Currents

.LIB EVAL.LIB
X1 3 2 7 4 6 UA741
R1 3 0 1MEG
V1 7 0 15
V2 0 4 15
V0 2 6 0
.END
