;
.lib eval.lib
xa 3 2 7 4 6 ua741
vp 7 0 +15
vn 4 0 -15
r1 2 5 1k
rs 9 10 300
d1 6 8 d1n4002
c1 5 9 .02u
rl 8 0 10k
vin 10 0 sin 0 2 1k
vref 3 0 1
.tran .1m 2m
.probe 
.end

