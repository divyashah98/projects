NON INVERTING AMPLIFIER

.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
V1 7 0 DC 15
V2 0 4 DC 15
Ra 2 0 1K
Rf 2 6 15K
Vs 3 0 SIN(0 100M 1K)
Rl 6 0 10k
.TRAN 500U 5M
.PROBE
.END
