Band Pass Filter
.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
Vp 7 0 15
Vn 0 4 15
Ra 1 5 1K
Ca 5 0 0.5U
Cb 5 3 0.5U
Rb 3 0 2K
Rc 5 6 1K
R1 2 0 1K
R2 6 2 1K
Vin 1 0 AC 100M
.AC DEC 20 10 10K
.PROBE
.END
