;
.lib eval.lib
xa 1 5 2 3 4 ua741
vp 2 0 dc 15
vn 3 0 dc -15
vs 7 0 sin(.001 1k)
r1 6 5 1k
rs 1 7 300
rl 4 0 10k
c1 6 0 .51u
d1 5 1 d1n4002
d2 1 5 d1n4002
.tran 0.1m 1k
.probe 
.end
