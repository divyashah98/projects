Positive Clamping Circuit

.LIB EVAL.LIB
.MODEL 1N4002 D
Xa 3 2 7 4 6 UA741
va 0 4 15
vb 7 0 15
VreF 3 0 30
Ra 2 9 100
Da 6 9 D1N4002
*.MODEL D1N4001 D (IS=18.8n RS=0 BV=400 IBV=5.00u CJO=30 M=0.333 N=2)
Rl 9 0 10K
Ca 9 1 100U IC 35
Vin 1 0 SIN(0 20 2k)
.TRAN 0.1m 10M 
.PROBE
.END
