Chopper
.lib nom.lib
Vdc 1 0 12
Jfet1 1 2 3 J2N3819
Vs1 2 0 pulse(0 -15 0 0.1n 0.1n 10u 20u)
D1 0 3 D1N4002
L1 3 4 16m
C1 4 0 100u
R1 4 0 100k
.probe
.tran 10u 200u
.end

