3_2
.LIB EVAL.LIB
Xa 3 2 7 4 6 UA741
D1 6 9 D1N4002
D2 0 6 D1N4002
Vp 7 0 15
Vn 0 4 15
Ra 3 1 300
Vin 1 0 SIN(0 5 1k)
Rb 2 9 1K
Rl 9 0 10K
Cl 9 0 0.2U
.TRAN 100u 5M
.PROBE
.END
