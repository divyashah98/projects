library verilog;
use verilog.vl_types.all;
entity prog_sqr_wav_gen_tb is
end prog_sqr_wav_gen_tb;
